----------------------------------------------------------------------------------
-- Company: UERGS
-- Disciplina: Organizacao de computadores
-- Profa.: Debora Matos
-- Baseado na estrutura de memoria de: Newton Jr
-- Trabalho de: Ismael Soller Vianna
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.NUMERIC_STD.ALL;
library mito;
use mito.mito_pkg.all;

entity memory is
	port(		
        clk                 : in  std_logic;
        escrita             : in  std_logic;                     -- habilita escrita em 1
        rst                 : in  std_logic;        
        entrada_memoria     : in  std_logic_vector(31 downto 0); -- dado a ser inserido na memoria
        endereco_memoria    : in  std_logic_vector(8  downto 0); -- endere�o a ser lido ou gravado
        saida_memoria       : out std_logic_vector(31 downto 0)
        );        
end memory;

architecture rtl of memory is

	-- 128 words of 4 bytes (32 bits)
	subtype palavra is std_logic_vector(7 downto 0);
	type memory is array (0 to 511) of palavra;
	signal mem : memory;
	
begin 

process(clk, escrita, endereco_memoria, rst)	
begin	
            if(rst = '1') then     
                mem(0)    <= "00101100";
                mem(1)    <= "00000001";
                mem(2)    <= "00000000";
                mem(3)    <= "00000101";
                mem(4)    <= "01111100";
                mem(5)    <= "00100010";
                mem(6)    <= "00000000";
                mem(7)    <= "10011111";
                mem(8)    <= "00011000";
                mem(9)    <= "00000000";
                mem(10)    <= "00000000";
                mem(11)    <= "00000000";
                mem(12)    <= "00001000";
                mem(13)    <= "00100010";
                mem(14)    <= "00000000";
                mem(15)    <= "00000001";
                mem(16)    <= "00101100";
                mem(17)    <= "00000101";
                mem(18)    <= "00000000";
                mem(19)    <= "00000011";
                mem(20)    <= "00100100";
                mem(21)    <= "00100100";
                mem(22)    <= "00011000";
                mem(23)    <= "00000001";
                mem(24)    <= "00011000";
                mem(25)    <= "00000000";
                mem(26)    <= "00000000";
                mem(27)    <= "00000000";
                mem(28)    <= "00011000";
                mem(29)    <= "00000000";
                mem(30)    <= "00000000";
                mem(31)    <= "00000000";
                mem(32)    <= "00101100";
                mem(33)    <= "00000010";
                mem(34)    <= "00000000";
                mem(35)    <= "00000111";
                mem(36)    <= "01101000";
                mem(37)    <= "01000001";
                mem(38)    <= "00000000";
                mem(39)    <= "00110000";
                mem(40)<= "00011000";
                mem(41)<= "00000000";
                mem(42)<= "00000000";
                mem(43)<= "00000000";
                mem(44)<= "00101100";
                mem(45)<= "00000010";
                mem(46)<= "00000000";
                mem(47)<= "00001010";
                mem(48)<= "00101100";
                mem(49)<= "00000001";
                mem(50)<= "00000000";
                mem(51)<= "00001011";
                mem(52)<= "00011000";
                mem(53)<= "00000000";
                mem(54)<= "00000000";
                mem(55)<= "00000000";
                mem(56)<= "00000000";
                mem(57)<= "00000000";
                mem(58)<= "00000000";
                mem(59)<= "00000000";
                mem(60)<= "00000000";
                mem(61)<= "00000000";
                mem(62)<= "00000000";
                mem(63)<= "00000000";
                mem(64)<= "00000000";
                mem(65)<= "00000000";
                mem(66)<= "00000000";
                mem(67)<= "00000000";
                mem(68)<= "00000000";
                mem(69)<= "00000000";
                mem(70)<= "00000000";
                mem(71)<= "00000000";
                mem(72)<= "00000000";
                mem(73)<= "00000000";
                mem(74)<= "00000000";
                mem(75)<= "00000000";
                mem(76)<= "00000000";
                mem(77)<= "00000000";
                mem(78)<= "00000000";
                mem(79)<= "00000000";
                mem(80)<= "00000000";
                mem(81)<= "00000000";
                mem(82)<= "00000000";
                mem(83)<= "00000000";
                mem(84)<= "00000000";
                mem(85)<= "00000000";
                mem(86)<= "00000000";
                mem(87)<= "00000000";
                mem(88)<= "00000000";
                mem(89)<= "00000000";
                mem(90)<= "00000000";
                mem(91)<= "00000000";
                mem(92)   <= "00000000";
                mem(93)   <= "00000000";
                mem(94)   <= "00000000";
                mem(95)   <= "00000000";
                mem(96)   <= "00000000";
                mem(97)   <= "00000000";
                mem(98)   <= "00000000";
                mem(99)   <= "00000000";
                mem(100)  <= "00000000"; 
                mem(101)  <= "00000000";
                mem(102)  <= "00000000"; 
                mem(103)  <= "00000000";
                mem(104)  <= "00000000";
                mem(105)  <= "00000000";
                mem(106)  <= "00000000";
                mem(107)  <= "00000000";
                mem(108)  <= "00000000";
                mem(109)  <= "00000000";
                mem(110)  <= "00000000";
                mem(111)  <= "00000000";
                mem(112)  <= "00000000";
                mem(113)  <= "00000000";
                mem(114)  <= "00000000";
                mem(115)  <= "00000000";
                mem(116)  <= "00000000";
                mem(117)  <= "00000000";
                mem(118)  <= "00000000";
                mem(119)  <= "00000000";
                mem(120)  <= "00000000";
                mem(121)  <= "00000000";
                mem(122)  <= "00000000";
                mem(123)  <= "00000000";
                mem(124)  <= "00000000";
                mem(125)  <= "00000000";
                mem(126)  <= "00000000";
                mem(127)  <= "00000000";
                mem(128)  <= "00000000";
                mem(129)  <= "00000000"; 
                mem(130)  <= "00000000"; 
                mem(131)  <= "00000000";
                mem(132)  <= "00000000";
                mem(133)  <= "00000000";
                mem(134)  <= "00000000";
                mem(135)  <= "00000000";
                mem(136)  <= "00000000";
                mem(137)  <= "00000000";
                mem(138)  <= "00000000";
                mem(139)  <= "00000000";
                mem(140)  <= "00000000";
                mem(141)  <= "00000000";
                mem(142)  <= "00000000";
                mem(143)  <= "00000000";
                mem(144)  <= "00000000";
                mem(145)  <= "00000000";
                mem(146)  <= "00000000";
                mem(147)  <= "00000000";
                mem(148)  <= "00000000";
                mem(149)  <= "00000000";
                mem(150)  <= "00000000";
                mem(151)  <= "00000000";
                mem(152)  <= "00000000";
                mem(153)  <= "00000000";
                mem(154)  <= "00000000";
                mem(155)  <= "00000000";
                mem(156)  <= "00000000";
                mem(157)  <= "00000000";
                mem(158)  <= "00000000";
                mem(159)  <= "00000000";
                mem(160)  <= "00000000";
                mem(161)  <= "00000000";
                mem(162)  <= "00000000";
                mem(163)  <= "00000000";
                mem(164)  <= "00000000";
                mem(165)  <= "00000000";
                mem(166)  <= "00000000";
                mem(167)  <= "00000000";
                mem(168)  <= "00000000";
                mem(169)  <= "00000000";
                mem(170)  <= "00000000";
                mem(171)  <= "00000000";
                mem(172)  <= "00000000";
                mem(173)  <= "00000000";
                mem(174)  <= "00000000";
                mem(175)  <= "00000000";
                mem(176)  <= "00000000";
                mem(177)  <= "00000000";
                mem(178)  <= "00000000";
                mem(179)  <= "00000000";
                mem(180)  <= "00000000";
                mem(181)  <= "00000000";
                mem(182)  <= "00000000";
                mem(183)  <= "00000000";
                mem(184)  <= "00000000";
                mem(185)  <= "00000000";
                mem(186)  <= "00000000";
                mem(187)  <= "00000000";
                mem(188)  <= "00000000";
                mem(189)  <= "00000000";
                mem(190)  <= "00000000";
                mem(191)  <= "00000000";
                mem(192)  <= "00000000";
                mem(193)  <= "00000000";
                mem(194)  <= "00000000";
                mem(195)  <= "00000000";
                mem(196)  <= "00000000";
                mem(197)  <= "00000000";
                mem(198)  <= "00000000";
                mem(199)  <= "00000000";
                mem(200)  <= "00000000";
                mem(201)  <= "00000000";
                mem(202)  <= "00000000";
                mem(203)  <= "00000000";
                mem(204)  <= "00000000";
                mem(205)  <= "00000000";
                mem(206)  <= "00000000";
                mem(207)  <= "00000000";
                mem(208)  <= "00000000";
                mem(209)  <= "00000000";
                mem(210)  <= "00000000";
                mem(211)  <= "00000000";
                mem(212)  <= "00000000";
                mem(213)  <= "00000000";
                mem(214)  <= "00000000";
                mem(215)  <= "00000000";
                mem(216)  <= "00000000";
                mem(217)  <= "00000000";
                mem(218)  <= "00000000";
                mem(219)  <= "00000000";
                mem(220)  <= "00000000";
                mem(221)  <= "00000000";
                mem(222)  <= "00000000";
                mem(223)  <= "00000000";
                mem(224)  <= "00000000";
                mem(225)  <= "00000000";
                mem(226)  <= "00000000";
                mem(227)  <= "00000000";
                mem(228)  <= "00000000";
                mem(229)  <= "00000000";
                mem(230)  <= "00000000";
                mem(231)  <= "00000000";
                mem(232)  <= "00000000";
                mem(233)  <= "00000000";
                mem(234)  <= "00000000";
                mem(235)  <= "00000000";
                mem(236)  <= "00000000";
                mem(237)  <= "00000000";
                mem(238)  <= "00000000";
                mem(239)  <= "00000000";
                mem(240)  <= "00000000";
                mem(241)  <= "00000000";
                mem(242)  <= "00000000";
                mem(243)  <= "00000000";
                mem(244)  <= "00000000";
                mem(245)  <= "00000000";
                mem(246)  <= "00000000";
                mem(247)  <= "00000000";
                mem(248)  <= "00000000";
                mem(249)  <= "00000000";
                mem(250)  <= "00000000";
                mem(251)  <= "00000000";
                mem(252)  <= "00000000";
                mem(253)  <= "00000000";
                mem(254)  <= "00000000";
                mem(255)  <= "00000000";
                mem(256)  <= "00000000";
                mem(257)  <= "00000000";
                mem(258)  <= "00000000";
                mem(259)  <= "00000000";
                mem(260)  <= "00000000";
                mem(261)  <= "00000000";
                mem(262)  <= "00000000";
                mem(263)  <= "00000000";
                mem(264)  <= "00000000";
                mem(265)  <= "00000000";
                mem(266)  <= "00000000";
                mem(267)  <= "00000000";
                mem(268)  <= "00000000";
                mem(269)  <= "00000000";
                mem(270)  <= "00000000";
                mem(271)  <= "00000000";
                mem(272)  <= "00000000";
                mem(273)  <= "00000000";
                mem(274)  <= "00000000";
                mem(275)  <= "00000000";
                mem(276)  <= "00000000";
                mem(277)  <= "00000000";
                mem(278)  <= "00000000";
                mem(279)  <= "00000000";
                mem(280)  <= "00000000";
                mem(281)  <= "00000000";
                mem(282)  <= "00000000";
                mem(283)  <= "00000000";
                mem(284)  <= "00000000";
                mem(285)  <= "00000000";
                mem(286)  <= "00000000";
                mem(287)  <= "00000000";
                mem(288)  <= "00000000";
                mem(289)  <= "00000000";
                mem(290)  <= "00000000";
                mem(291)  <= "00000000";
                mem(292)  <= "00000000";
                mem(293)  <= "00000000";
                mem(294)  <= "00000000";
                mem(295)  <= "00000000";
                mem(296)  <= "00000000";
                mem(297)  <= "00000000";
                mem(298)  <= "00000000";
                mem(299)  <= "00000000";
                mem(300)  <= "00000000";
                mem(301)  <= "00000000";
                mem(302)  <= "00000000";
                mem(303)  <= "00000000";
                mem(304)  <= "00000000";
                mem(305)  <= "00000000";
                mem(306)  <= "00000000";
                mem(307)  <= "00000000";
                mem(308)  <= "00000000";
                mem(309)  <= "00000000";
                mem(310)  <= "00000000";
                mem(311)  <= "00000000";
                mem(312)  <= "00000000";
                mem(313)  <= "00000000";
                mem(314)  <= "00000000";
                mem(315)  <= "00000000";
                mem(316)  <= "00000000";
                mem(317)  <= "00000000";
                mem(318)  <= "00000000";
                mem(319)  <= "00000000";
                mem(320)  <= "00000000";
                mem(321)  <= "00000000";
                mem(322)  <= "00000000";
                mem(323)  <= "00000000";
                mem(324)  <= "00000000";
                mem(325)  <= "00000000";
                mem(326)  <= "00000000";
                mem(327)  <= "00000000";
                mem(328)  <= "00000000";
                mem(329)  <= "00000000"; 
                mem(330)  <= "00000000"; 
                mem(331)  <= "00000000";
                mem(332)  <= "00000000";
                mem(333)  <= "00000000";
                mem(334)  <= "00000000";
                mem(335)  <= "00000000";
                mem(336)  <= "00000000";
                mem(337)  <= "00000000";
                mem(338)  <= "00000000";
                mem(339)  <= "00000000";
                mem(340)  <= "00000000";
                mem(341)  <= "00000000";
                mem(342)  <= "00000000";
                mem(343)  <= "00000000";
                mem(344)  <= "00000000";
                mem(345)  <= "00000000";
                mem(346)  <= "00000000";
                mem(347)  <= "00000000";
                mem(348)  <= "00000000";
                mem(349)  <= "00000000";
                mem(350)  <= "00000000";
                mem(351)  <= "00000000";
                mem(352)  <= "00000000";
                mem(353)  <= "00000000";
                mem(354)  <= "00000000";
                mem(355)  <= "00000000";
                mem(356)  <= "00000000";
                mem(357)  <= "00000000";
                mem(358)  <= "00000000";
                mem(359)  <= "00000000";
                mem(360)  <= "00000000";
                mem(361)  <= "00000000";
                mem(362)  <= "00000000";
                mem(363)  <= "00000000";
                mem(364)  <= "00000000";
                mem(365)  <= "00000000";
                mem(366)  <= "00000000";
                mem(367)  <= "00000000";
                mem(368)  <= "00000000";
                mem(369)  <= "00000000";
                mem(370)  <= "00000000";
                mem(371)  <= "00000000";
                mem(372)  <= "00000000";
                mem(373)  <= "00000000";
                mem(374)  <= "00000000";
                mem(375)  <= "00000000";
                mem(376)  <= "00000000";
                mem(377)  <= "00000000";
                mem(378)  <= "00000000";
                mem(379)  <= "00000000";
                mem(380)  <= "00000000";
                mem(381)  <= "00000000";
                mem(382)  <= "00000000";
                mem(383)  <= "00000000";
                mem(384)  <= "00000000";
                mem(385)  <= "00000000";
                mem(386)  <= "00000000";
                mem(387)  <= "00000000";
                mem(388)  <= "00000000";
                mem(389)  <= "00000000";
                mem(390)  <= "00000000";
                mem(391)  <= "00000000";
                mem(392)  <= "00000000";
                mem(393)  <= "00000000";
                mem(394)  <= "00000000";
                mem(395)  <= "00000000";
                mem(396)  <= "00000000";
                mem(397)  <= "00000000";
                mem(398)  <= "00000000";
                mem(399)  <= "00000000";
                mem(400)  <= "00000000";
                mem(401)  <= "00000000";
                mem(402)  <= "00000000";
                mem(403)  <= "00000000";
                mem(404)  <= "00000000";
                mem(405)  <= "00000000";
                mem(406)  <= "00000000";
                mem(407)  <= "00000000";
                mem(408)  <= "00000000";
                mem(409)  <= "00000000";
                mem(410)  <= "00000000";
                mem(411)  <= "00000000";
                mem(412)  <= "00000000";
                mem(413)  <= "00000000";
                mem(414)  <= "00000000";
                mem(415)  <= "00000000";
                mem(416)  <= "00000000";
                mem(417)  <= "00000000";
                mem(418)  <= "00000000";
                mem(419)  <= "00000000";
                mem(420)  <= "00000000";
                mem(421)  <= "00000000";
                mem(422)  <= "00000000";
                mem(423)  <= "00000000";
                mem(424)  <= "00000000";
                mem(425)  <= "00000000";
                mem(426)  <= "00000000";
                mem(427)  <= "00000000";
                mem(428)  <= "00000000";
                mem(429)  <= "00000000";
                mem(430)  <= "00000000";
                mem(431)  <= "00000000";
                mem(432)  <= "00000000";
                mem(433)  <= "00000000";
                mem(434)  <= "00000000";
                mem(435)  <= "00000000";
                mem(436)  <= "00000000";
                mem(437)  <= "00000000";
                mem(438)  <= "00000000";
                mem(439)  <= "00000000";
                mem(440)  <= "00000000";
                mem(441)  <= "00000000";
                mem(442)  <= "00000000";
                mem(443)  <= "00000000";
                mem(444)  <= "00000000";
                mem(445)  <= "00000000";
                mem(446)  <= "00000000";
                mem(447)  <= "00000000";
                mem(448)  <= "00000000";
                mem(449)  <= "00000000";
                mem(450)  <= "00000000";
                mem(451)  <= "00000000";
                mem(452)  <= "00000000";
                mem(453)  <= "00000000";
                mem(454)  <= "00000000";
                mem(455)  <= "00000000";
                mem(456)  <= "00000000";
                mem(457)  <= "00000000";
                mem(458)  <= "00000000";
                mem(459)  <= "00000000";
                mem(460)  <= "00000000";
                mem(461)  <= "00000000";
                mem(462)  <= "00000000";
                mem(463)  <= "00000000";
                mem(464)  <= "00000000";
                mem(465)  <= "00000000";
                mem(466)  <= "00000000";
                mem(467)  <= "00000000";
                mem(468)  <= "00000000";
                mem(469)  <= "00000000";
                mem(470)  <= "00000000";
                mem(471)  <= "00000000";
                mem(472)  <= "00000000";
                mem(473)  <= "00000000";
                mem(474)  <= "00000000";
                mem(475)  <= "00000000";
                mem(476)  <= "00000000";
                mem(477)  <= "00000000";
                mem(478)  <= "00000000";
                mem(479)  <= "00000000";
                mem(480)  <= "00000000";
                mem(481)  <= "00000000";
                mem(482)  <= "00000000";
                mem(483)  <= "00000000";
                mem(484)  <= "00000000";
                mem(485)  <= "00000000";
                mem(486)  <= "00000000";
                mem(487)  <= "00000000";
                mem(488)  <= "00000000";
                mem(489)  <= "00000000";
                mem(490)  <= "00000000";
                mem(491)  <= "00000000";
                mem(492)  <= "00000000";
                mem(493)  <= "00000000";
                mem(494)  <= "00000000";
                mem(495)  <= "00000000";
                mem(496)  <= "00000000";
                mem(497)  <= "00000000";
                mem(498)  <= "00000000";
                mem(499)  <= "00000000";
                mem(500)  <= "00000000";
                mem(501)  <= "00000000";
                mem(502)  <= "00000000";
                mem(503)  <= "00000000";
                mem(504)  <= "00000000";
                mem(505)  <= "00000000";
                mem(506)  <= "00000000";
                mem(507)  <= "00000000";
                mem(508)  <= "00000000";
                mem(509)  <= "00000000";
                mem(510)  <= "00000000";
                mem(511)  <= "00000000";
        else
            -- lendo da memoria
            if (escrita = '0') then                     
                    saida_memoria(31 downto 24) <= mem(to_integer(unsigned(endereco_memoria)));
                    saida_memoria(23 downto 16) <= mem(to_integer(unsigned(endereco_memoria+1)));
                    saida_memoria(15 downto  8) <= mem(to_integer(unsigned(endereco_memoria+2)));
                    saida_memoria( 7 downto  0) <= mem(to_integer(unsigned(endereco_memoria+3)));
                    
            -- escrevendo na memoria
            elsif (escrita = '1') then 		
                mem(to_integer(unsigned(endereco_memoria)))   <= entrada_memoria(31 downto 24);			
                mem(to_integer(unsigned(endereco_memoria+1))) <= entrada_memoria(23 downto 16);
                mem(to_integer(unsigned(endereco_memoria+2))) <= entrada_memoria(15 downto  8);
                mem(to_integer(unsigned(endereco_memoria+3))) <= entrada_memoria( 7 downto  0);
                
            end if;
        end if;		    					
end process;

end rtl;
